// Design a multiplier circuit that does multiplication of two 16-bit inputs by repeatative addition.
