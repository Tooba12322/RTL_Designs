module comp_2b
