// From input code, generate 7 segment code and print its respective ASCII value
