//16-bit ripple carry adder - structural modeling

module 


endmodule
