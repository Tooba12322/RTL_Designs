// Waveform : 
//mode-0 (cpol=0,cpha=0) https://www.edaplayground.com/w/x/Cid
//mode-1 (cpol=0,cpha=1) https://www.edaplayground.com/w/x/Fp5
//mode-2 (cpol=1,cpha=0) https://www.edaplayground.com/w/x/JtW
//mode-3 (cpol=1,cpha=1) https://www.edaplayground.com/w/x/RgE

`timescale 1ns/1ps
module spi_s_tb();
 
  logic done,miso;
  logic [7:0] dout;
  logic mosi,rst,cpha,cpol,sclk,ready; // no system clk, it runs on sclk generated by master
  logic [7:0] din;
  
  spi_s DUT(.*);
    
 initial
  begin
    $dumpfile("spi_s.vcd");
    $dumpvars(0,spi_s_tb);
    
    rst      = '0;
    mosi     = '0;
    din      = '0;
    cpol     = '1;
    cpha     = '1;
    ready    = '1;
    sclk     = '0;
    
    #7  rst = '1;

    #7 din = 8'hA1;
    ready = (!done) ? '0 : '1;
    

    for (int i=0;i<20;i++) begin
      mosi = $random%6 || $random%3;
      sclk = !sclk;
      #550;
    end
   #10 $finish;
  end
 
endmodule
