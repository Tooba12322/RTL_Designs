// Design a gray code counter that generates all 4-bit and 3-bit gray counts.
// n-bit and (n-1) bit gray counter, the (n-1)-bit Gray code is simply generated 
// by doing an exclusive-or operation on the two MSBs of the n-bit Gray code
// to generate the MSB for the (n-1)-bit Gray code.
// This is combined with the (n-2) LSBs of the n-bit Gray code counter to form the (n-1)-bit Gray code counter.
