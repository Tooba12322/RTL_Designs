// Command interface design, using it inside a module
