// Design a circuit that detects the sequence "0110" without overlapping, from continuous bit stream.
