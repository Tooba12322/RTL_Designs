// Variable swapping using blocking and non-blocking statements
