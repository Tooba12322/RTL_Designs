// Async mod-10 counter
