//Design a Moore FSM to control a traffic light system. 
//The FSM should have three states corresponding to the traffic light colors: Red, Green, and Yellow. 
//The traffic light should cycle through these states in the order Red → Green → Yellow → Red, with a fixed time duration for each color. 
//The FSM should have a clock input for timing and a reset input to restart the cycle. The output should indicate the current color of the traffic light.
