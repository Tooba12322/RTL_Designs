// Design a sequence detector to detect "101010" in overlapping fashion using Mealey FSM
