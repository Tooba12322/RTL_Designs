// Design a circiut whose output is the GCD (Greatest Common Deviser) of two integers, using continuous subtraction algorithm
