module D_latch()

endmodule

module SR_latch()

endmodule
