// Design a circuit that identifies parity of input bit steam,even=1,odd=0
