// Design a UART system with both transmission and reception functionality ,
// use FIFOs to transmit/recieve data from/to fast running CPU 
