// Implement an 8-bit counter
  // - Resets to 0
  // - Increments by 1 every cycle
  // - Takes the load value if load_i is seen
  // - Starts to count down after overflow, otherwise count up
  
