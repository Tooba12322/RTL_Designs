// Design a circuit that detects three or more consequtive 1's in the continuous bit stream.
