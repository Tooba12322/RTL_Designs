// Debouncing circuit implementation usin delayed detection with delay equals to 2-3msec
