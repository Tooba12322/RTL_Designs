module D_latch_tb()

endmodule

module SR_latch_tb()

endmodule
