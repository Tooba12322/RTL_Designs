module LUT(F,a0, a1, a2, a3, clk, rst);
  logic F;
  logic a0, a1, a2, a3;
  logic clk;
  logic rst;
  logic RAM[15:0];
  
endmodule

